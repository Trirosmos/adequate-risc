module cpu(
	input clk
);

reg [27:0] pc;

wire advance_pc = pc + 1;



endmodule